// this is the top tesbench UVM file

`timescale 1ns/1ns

import uvm_pkg::*;
`include "uvm_macros.svh"

module top;







endmodule: top